module axi_slave(

	  input[31:0] M_AXI_GP0_araddr,
	  input[1:0] M_AXI_GP0_arburst,
	  input[3:0] M_AXI_GP0_arcache,
	  input[11:0] M_AXI_GP0_arid,
	  input[3:0] M_AXI_GP0_arlen,
	  input[1:0] M_AXI_GP0_arlock,
	  input[2:0] M_AXI_GP0_arprot,
	  input[3:0] M_AXI_GP0_arqos,
	  output M_AXI_GP0_arready,
	  input[2:0] M_AXI_GP0_arsize,
	  input M_AXI_GP0_arvalid,
	  input[31:0] M_AXI_GP0_awaddr,
	  input[1:0] M_AXI_GP0_awburst,
	  input[3:0] M_AXI_GP0_awcache,
	  input[11:0] M_AXI_GP0_awid,
	  input[3:0] M_AXI_GP0_awlen,
	  input[1:0] M_AXI_GP0_awlock,
	  input[2:0] M_AXI_GP0_awprot,
	  input[3:0] M_AXI_GP0_awqos,
	  output M_AXI_GP0_awready,
	  input[2:0] M_AXI_GP0_awsize,
	  input M_AXI_GP0_awvalid,
	  output [11:0] M_AXI_GP0_bid,
	  input M_AXI_GP0_bready,
	  output [1:0] M_AXI_GP0_bresp,
	  output M_AXI_GP0_bvalid,
	  output [31:0] M_AXI_GP0_rdata,
	  output [11:0] M_AXI_GP0_rid,
	  output M_AXI_GP0_rlast,
	  input M_AXI_GP0_rready,
	  output [1:0] M_AXI_GP0_rresp,
	  output M_AXI_GP0_rvalid,
	  input[31:0] M_AXI_GP0_wdata,
	  input[11:0] M_AXI_GP0_wid,
	  input M_AXI_GP0_wlast,
	  output M_AXI_GP0_wready,
	  input[3:0] M_AXI_GP0_wstrb,
	  input M_AXI_GP0_wvalid
	  );
  

endmodule // axi_slave